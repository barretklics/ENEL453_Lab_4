/*module FM_Modulator #(parameter int
							min_dist = 400,
							max_dist = 2000
							)
							
	(input logic [11:0] distance,
	output logic tuning_word
	);
	
	
	
	
	
	
	
	
	
	
	always_comb 
	begin
	
	
	
	
	
         
	end
	
	
	
	
	
	
endmodule*/