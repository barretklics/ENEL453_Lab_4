module debug_module
 #(parameter width=16)
	(output logic [width-1:0] debug_out
	);

	  
  assign debug_out = 16'b0101101001011010;
  
  endmodule